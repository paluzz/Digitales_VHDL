-- ej1: entradas A y B , si sel = 0 -> RES = A + B en magnitud (unsigned)
--                      si sel = 1 -> RES = A + B en CA2 (signed)

-- ej2: si sel1 = 0 -> comp = A si A > B
--      si sel2 = 1 -> comp = A si A < B

-- ej3: TOP level con dos comparadores y un sumador
--
architecture rtl of comp is
begin
end architecture;